`timescale 1ns / 100ps
//
//////////////////////////////////////////////////////////////////////////////////
//
//  Filename: tb_multicycle.sv
//
//  Author: Mike Wirthlin
//  
//////////////////////////////////////////////////////////////////////////////////

module tb_multicycle #(
    TEXT_ADDRESS = 32'h00200000,
    DATA_ADDRESS = 32'h00000000,
    string instruction_memory_filename = "simple_datapath_text.mem",
    string data_memory_filename = "simple_datapath_data.mem",
    int MAX_INSTRUCTION_COUNT = 2000
    ) ();

    import tb_riscv_pkg::*;

    // Testbench global signals
    logic clk, rst;
    // DUT input signals (used by DUT)
    logic [31:0] instruction;
    logic [31:0] dReadData;
    // // DUT output sigals (generated by DUT)
    logic [31:0] PC;
    logic [31:0] dWriteData, dAddress, WriteBackData;
    logic MemRead, MemWrite;

    // clock generation
    initial begin
        clk = 0;
        forever #5 clk <= ~clk; // 100MHz
    end

    // Instance Datapath module
    riscv_multicycle #(.INITIAL_PC(TEXT_ADDRESS))
    riscv_multicycle(.*);

    // Instance simulation model
    riscv_simple_datapath_model #(
        .TEXT_ADDRESS(TEXT_ADDRESS),
        .instruction_memory_filename(instruction_memory_filename),
        .data_memory_filename(data_memory_filename)
    ) riscv_model(
        // Testbench inputs
        .clk(clk), .rst(rst),
        // Control Signals to drive to DUT (for datapath lab)
        .PCSrc(), .loadPC(), .ALUSrc(), .RegWrite(), .MemtoReg(), .ALUCtrl(),
        // Memory interface signals
        .instruction(instruction), .dAddress(dAddress),
        .dWriteData(dWriteData), .dReadData(dReadData),
        // Signals to check
        // .Zero(Zero),
        .PC(PC), .WriteBackData(WriteBackData)
    );

    initial begin

        //shall print %t with scaled in ns (-9), with 2 precision digits, and would print the " ns" string
        $timeformat(-9, 0, " ns", 20);
        $display("*** Start of Simulation ***");

        // Initialize the inputs
        repeat(3) @(negedge clk);
        rst = 1;
        repeat(3) @(negedge clk);
        rst = 0;

        while(instruction != riscv_instr::EBREAK_INSTRUCTION) begin
            @(negedge clk);
            if (riscv_model.error != 0) begin
                $display("*** Simulation stopped due to error @ %0t *** ", $time);
                $finish;
            end
            if (riscv_model.instruction_count >= MAX_INSTRUCTION_COUNT) begin
                $display("*** Simulation stopped due to max instruction count (%0d) @ %0t *** ",
                    MAX_INSTRUCTION_COUNT, $time);
                $finish;
            end
        end

        $display("*** Simulation done @ %0t - %0d instructions *** ", $time, riscv_model.instruction_count);
        if (riscv_model.error == 0)
            $display("===== TEST PASSED =====");
        else
            $display("===== TEST FAILED =====");

        $finish;

    end  // end initial
    
endmodule

// This model simulates the datapath and generates the control signals for testing.
module riscv_simple_datapath_model #(
    string instruction_memory_filename,
    string data_memory_filename,
    logic [31:0] TEXT_ADDRESS = 32'h00200000,
    logic [31:0] DATA_ADDRESS = 32'h00000000,
    int MAX_TEXT_SIZE = 4096,
    int MAX_DATA_SIZE = 1024
    ) 
    (
        input logic clk,
        input logic rst,
        // Control signals for student datapath module
        output logic PCSrc,
        output logic loadPC,
        output logic ALUSrc,
        output logic RegWrite,
        output logic MemtoReg,
        output logic [3:0] ALUCtrl,
        // Memory interface signals to DUT
        output logic [31:0] instruction,
        output logic [31:0] dReadData,
        // Signals from DUT to check:
        input logic Zero,
        input [31:0] PC,
        input MemRead,
        input MemWrite,
        input [31:0] dWriteData,
        input [31:0] dAddress,
        input [31:0] WriteBackData
    );

    import tb_riscv_pkg::*;

    typedef enum { IF, ID, EX, MEM, WB } inst_stage_t;
    inst_stage_t current_stage;

    riscv_regfile regfile;
    riscv_instr cur_inst;
    riscv_simple_control riscv_ctrl;

    logic tb_alu_Zero;
    logic [31:0] tb_alu, readA, readB, b_operand, tb_writeBackData;
    logic [31:0] PC_i, dAddress_i, dWriteData_i, dReadData_i;
    logic MemRead_i, MemWrite_i;

     // Instruction Memory
    logic error = 0;
    int instruction_count = 0;
    logic initialized = 0;

    // Instruction Memory (don't print memory transactions for instruction memory)
    riscv_memory #(
        .MEMORY_FILENAME(instruction_memory_filename), .MEMORY_NAME(".text"),
        .MEMORY_WORDS(MAX_TEXT_SIZE), .MEMORY_OFFSET(TEXT_ADDRESS),
        .PRINT_MEMORY_TRANSACTIONS(0), .DEFAULT_MEMORY_VALUE(NOP_INSTRUCTION)
    ) instruction_memory(
        .clk(clk), .rst(rst),
        .read_en(1'b1), .write_en(1'b0), .address(PC_i),
        .write_data('0), .read_data(instruction)
    );

    // Data Memory
    assign dAddress_i = tb_alu;
    assign dWriteData_i = readB;
    riscv_memory #(
        .MEMORY_FILENAME(data_memory_filename), .MEMORY_NAME(".data"),
        .MEMORY_WORDS(MAX_DATA_SIZE), .MEMORY_OFFSET(DATA_ADDRESS),
        .PRINT_MEMORY_TRANSACTIONS(0), .DEFAULT_MEMORY_VALUE(32'h00000000)
    ) data_memory(
        .clk(clk), .rst(rst),
        .read_en(MemRead_i), .write_en(MemWrite_i), .address(dAddress_i),
        .write_data(dWriteData_i), .read_data(dReadData_i)
    );

    initial begin
        regfile = new();
    end

    assign dReadData = dReadData_i;
    always_ff @(posedge clk or posedge rst) begin
        if (rst) begin
            // Internal signals
            current_stage <= IF;
            // Control signals
            loadPC <= 0;
            PCSrc <= 0;
            ALUSrc <= 0;
            RegWrite <= 0;
            MemtoReg <= 0;
            ALUCtrl <= 0;
            error <= 0;
            PC_i <= TEXT_ADDRESS;
            if (!initialized)
                $display("[%0t] rst Asserted", $time);
            initialized <= 1;
        end else if (initialized === 1'b1) begin
            MemRead_i <= 0;
            MemWrite_i <= 0;
            // dReadData <= 32'hxxxxxxxx;
            case (current_stage)
                IF: begin // End of IF stage/start of ID stage
                    #1step;
                    current_stage <= ID;
                end
                ID: begin // End of ID stage
                    #1step;
                    current_stage <= EX;
                    riscv_ctrl = new(instruction);
                    readA = regfile.read_rs1_i(instruction);
                    readB = regfile.read_rs2_i(instruction);
                    b_operand = riscv_ctrl.b_operand(readB);
                end
                EX: begin // End of EX stage/start of MEM stage
                    #1step;
                    current_stage <= MEM;
                    // Read Memory if needed (this is the start of MEM)
                    if (riscv_ctrl.MemRead)
                        MemRead_i <= 1;
                    if (riscv_ctrl.MemWrite)
                        MemWrite_i <= 1;
                end
                MEM: begin // End of MEM stage/start of WB stage
                    #1step;
                    current_stage <= WB;
                    // Display valid read data only on MemRead (during WB stage)
                    // if (riscv_ctrl.MemRead)
                    //     dReadData <= dReadData_i;
                    // // Write Memory
                    // if (riscv_ctrl.MemWrite) begin
                    //     data_mem.write(tb_alu >> 2, readB);
                    // end
                end
                WB: begin
                    #1step;
                    // if (riscv_ctrl.MemRead)
                    //     dReadData <= dReadData_i;
                    current_stage <= IF;
                    instruction_count = instruction_count + 1;
                    if (RegWrite)
                        regfile.write_reg_i(instruction, tb_writeBackData);
                    if (PCSrc) PC_i = PC_i + cur_inst.imm_b();
                    else PC_i = PC_i + 4;
                    RegWrite = 0;
                    loadPC = 0;
                end
            endcase
        end
    end

    always_ff @(negedge clk) begin
        if (initialized === 1'b1 && rst == 0) begin
            case (current_stage)
                IF: begin // ID stage
                    $display("==========================");
                    $display("[%0t] IF:  PC=%08h ", $time, PC_i);
                    if (PC_i != PC || ^PC[0] === 1'bX) begin
                        $display("**** Error: PC=%h but expect %h at time %0t", PC, PC_i, $time);
                        error = 1;
                    end
                end
                ID: begin
                    cur_inst = new(instruction);
                    $display("[%0t] ID:  INST=%08x %s", $time, cur_inst.u, cur_inst.inst_str());
                    riscv_ctrl = new(instruction);
                    ALUCtrl = riscv_ctrl.ALUCtrl;
                    ALUSrc = riscv_ctrl.ALUSrc;
                    // No checking here
                end
                EX: begin
                    tb_alu = riscv_alu::exec(riscv_alu::aluop_t'(ALUCtrl), readA, b_operand);
                    tb_alu_Zero = (tb_alu == 0);
                    $display("[%0t] EX:  dAddress=%08h zero=%b", $time, tb_alu, tb_alu_Zero);
                    // dAddress is the address to the data memory (or ALU result output)
                    if (tb_alu != dAddress || ^dAddress[0] === 1'bX) begin
                        $display("*** Error: dAddress=%h but expect %h at time %0t", dAddress, tb_alu, $time);
                        error = 1;
                        // error();
                    end else
                    if (tb_alu_Zero != Zero || Zero == 1'bX) begin
                        $display("*** Error: Zero=%h but expect %h at time %0t", Zero,
                        tb_alu_Zero, $time);
                        error = 1;
                        // error();
                    end
                end
                MEM: begin
                    // The write data is just the readB value from the register file
                    $write("[%0t] MEM: dWriteData=%08h", $time, readB);
                    if (riscv_ctrl.MemRead)
                        $display(" (MemRead)");
                    else if (riscv_ctrl.MemWrite)
                        $display(" (MemWrite)");
                    else
                        $display("");
                end
                WB: begin
                    loadPC = 1;        // prepare for next IF stage (this is put in WB instead of IF so the first cycle works correctly)
                    current_stage = WB;
                    RegWrite = riscv_ctrl.RegWrite;
                    MemtoReg = riscv_ctrl.MemtoReg;
                    tb_writeBackData = MemtoReg ? dReadData : tb_alu;
                    PCSrc = tb_alu_Zero & riscv_ctrl.branch;
                    $display("[%0t] WB:  WriteBackData=%08h", $time, tb_writeBackData);
                    // Check WriteBackData
                    if (RegWrite && (WriteBackData != tb_writeBackData || ^WriteBackData[0] === 1'bX)) begin
                        $display("*** Error: WriteBackData=%h but expect %h at time %0t", WriteBackData,
                        tb_writeBackData, $time);
                        error = 1;
                    end
                end
            endcase
        end
    end

endmodule