`timescale 1ns / 100ps
//
//////////////////////////////////////////////////////////////////////////////////
//
//  Filename: tb_simple_datapath.v
//
//  Author: Mike Wirthlin
//  
//////////////////////////////////////////////////////////////////////////////////

module tb_simple_datapath #(
    TB_INITIAL_PC = 32'h00200000,
    parameter instruction_memory_filename = "simple_datapath_text.mem",
    parameter data_memory_filename = "simple_datapath_data.mem",
    int MAX_TEXT_SIZE = 2048,
    int MAX_DATA_SIZE = 64
    ) ();

    import tb_riscv_pkg::*;

    // DUT input signals (used by DUT)
    logic clk, rst;
    logic PCSrc, loadPC, ALUSrc, RegWrite, MemtoReg; 
    logic [3:0] ALUCtrl;
    logic [31:0] instruction;
    logic [31:0] dReadData;
    // DUT output sigals (generated by DUT)
    logic [31:0] PC;
    logic [31:0] dWriteData, dAddress, WriteBackData;
    logic Zero;
    // Testbench signals
    riscv_instr cur_inst;
    riscv_simple_control riscv_ctrl;
    logic [31:0] tb_alu;
    logic tb_alu_Zero;
    logic [31:0] tb_readA, tb_readB, tb_b_operand, tb_writeData;
    logic [31:0] tb_PC;
    // integer i;
    // Simulation models
    riscv_regfile regfile;
    riscv_mem inst_mem;
    riscv_mem data_mem;

    typedef enum { IF, ID, EX, MEM, WB } inst_stage_t;
    inst_stage_t current_stage;

    // clock generation
    initial begin
        clk = 0;
        forever #5 clk <= ~clk; // 100MHz cl    typedef enum { IF, ID, EX, MEM, WB } inst_stage_t;
    end

    // Instance Datapath module
    riscv_simple_datapath #(.INITIAL_PC(TB_INITIAL_PC)) datapath(.*);

    task init_control();
        // Initializes all of the control signals to zero
        loadPC = 0;
        PCSrc = 0;
        ALUSrc = 0;
        RegWrite = 0;
        ALUCtrl = 0;
        MemtoReg = 0;
        instruction = '0;
        // Testbench signals
        tb_alu = 0;
        tb_alu_Zero = 0;
        tb_readA = 0;
        tb_readB = 0;
        tb_b_operand = 0;
        tb_writeData = 0;
    endtask

    task error();
        // Provide some delay after error so that you don't have to look at end of waveform
        #10 clk = 0;
        //$error;
        $finish;
    endtask;

    // assume currently at negative edge of clock
    task execute_instruction;
        begin
            if_stage();
            id_stage();
            ex_stage();
            mem_stage();
            wb_stage();
        end
    endtask

    // Each of the 'stage' tasks assume that they start at the negative edge of the
    // current stage and end at the negative edge of next stage
    // State at the end of the stage is updated on the positive edge of the clock 
    //  (in the middle of the task)
    // Stimulus is set on the negative edges and results are checked on the negative edges.

    // if_stage: (begin on neg edge of 'if' stage and end on neg edge of next 'id' stage)
    //  start edge: new PC, middle: initiale instruction read, end edge: new instruction
    // - clk action: update the PC for the new instruction
    // - neg edge check: PC is correct
    // - neg edge action: clear loadPC (so PC is not updated on next clock cycle)
    task automatic if_stage;
        current_stage = IF;
        $display("==========================");
        $display("[%0t] IF:  PC=%08h ", $time, tb_PC);
        @(negedge clk);
        if (tb_PC != PC || ^PC[0] === 1'bX) begin
            $display("*** Error: PC=%h but expect %h at time %0t", PC, tb_PC, $time);
            error();
        end
        @(posedge clk);
        #1step;
        // Read the current instruction
        instruction = inst_mem.read((tb_PC - TB_INITIAL_PC) >> 2);
        cur_inst = new(instruction);
    endtask

    // id_stage: (begin on neg edge of previous 'if' stage)
    // - clk action: read instruction from instruction memory
    // - neg edge action: set ALUCtrl and ALUSrc (i.e., decoding instruction)
    // - neg edge check: No checks since TB owns the instruction memory
    task id_stage;
        current_stage = ID;
        $display("[%0t] ID:  INST=%08x %s", $time, cur_inst.u, cur_inst.inst_str());
        @(negedge clk);
        riscv_ctrl = new(instruction);
        ALUCtrl = riscv_ctrl.ALUCtrl;
        ALUSrc = riscv_ctrl.ALUSrc;
        @(posedge clk);
        #1step;
        // Read the register file
        tb_readA = regfile.read_rs1_i(instruction);
        tb_readB = regfile.read_rs2_i(instruction);
        tb_b_operand = riscv_ctrl.b_operand(tb_readB);
    endtask

    // ex_stage: (begin on neg edge of previous 'id' stage)
    // - clk action: read the register file from the decoded instruction, compute updated tb ALU values
    // - neg edge check: check tb_alu and tb_alu_Zero against dAddress and Zero
    task ex_stage;
        current_stage = EX;
        tb_alu = riscv_alu::exec(riscv_alu::aluop_t'(ALUCtrl), tb_readA, tb_b_operand);
        tb_alu_Zero = (tb_alu == 0);
        $display("[%0t] EX:  dAddress=%08h zero=%b", $time, tb_alu, tb_alu_Zero);
        @(negedge clk);
        if (instruction != riscv_instr::EBREAK_INSTRUCTION) begin // ignore ebreak checks
            // dAddress is the address to the data memory (or ALU result output)
            if (tb_alu != dAddress || ^dAddress[0] === 1'bX) begin
                $display("*** Error: dAddress=%h but expect %h at time %0t", dAddress, tb_alu, $time);
                error();
            end else
            if (tb_alu_Zero != Zero || Zero == 1'bX) begin
                $display("*** Error: Zero=%h but expect %h at time %0t", Zero,
                tb_alu_Zero, $time);
                error();
            end
        end
        @(posedge clk);
        #1step;
    endtask

    // mem_stage: (begin on neg edge of previous 'ex' stage)
    // - clk action: read the register file from the decoded instruction, compute updated tb ALU values
    // - neg edge check: check tb_alu and tb_alu_Zero against dAddress and Zero


    task mem_stage;
        current_stage = MEM;
        // The write data is just the readB value from the register file
        $write("[%0t] MEM: dWriteData=%08h", $time, tb_readB);
        if (riscv_ctrl.MemRead)
            $display(" (MemRead)");
        else if (riscv_ctrl.MemWrite)
            $display(" (MemWrite)");
        else
            $display("");
        @(negedge clk);
        // Testbench provides the MemRead and MemWrite signals (but they don't go to the DUT)

        // Does the data to write match?
        if (riscv_ctrl.MemWrite && (dWriteData != tb_readB || ^dWriteData[0] === 1'bX ) ) begin
            $display("*** Error: dWriteData=%h but expect %h at time %0t", dWriteData,
            tb_readB, $time);
            error();
        end else
        // Don't need to check address since that would have been checked in EX stage

        @(posedge clk);
        #1step;
        // Write Memory
        if (riscv_ctrl.MemWrite) begin
            data_mem.write(tb_alu >> 2, tb_readB);
        end
        // Read Memory if needed
        if (riscv_ctrl.MemRead) begin
            dReadData = data_mem.read(tb_alu >> 2);
            // $display("[%0t] mem read %08h %0x %0x", $time, dReadData, tb_alu >> 2, tb_alu);
        end
        else
            dReadData = 32'hxxxxxxxx;
    endtask

    // activate: set pcsrc and regwrite. Provide read result
    // check: writebackdata
    task wb_stage;
        loadPC = 1;        // prepare for next IF stage (this is put in WB instead of IF so the first cycle works correctly)
        current_stage = WB;
        RegWrite = riscv_ctrl.RegWrite;
        MemtoReg = riscv_ctrl.MemtoReg;
        tb_writeData = MemtoReg ? dReadData : tb_alu;
        PCSrc = tb_alu_Zero & riscv_ctrl.branch;
        $display("[%0t] WB:  WriteBackData=%08h", $time, tb_writeData);
        @(negedge clk);
        // Check WriteBackData
        if (instruction != riscv_instr::EBREAK_INSTRUCTION && 
            RegWrite && (WriteBackData != tb_writeData || ^WriteBackData[0] === 1'bX)) begin
            $display("*** Error: WriteBackData=%h but expect %h at time %0t", WriteBackData,
            tb_writeData, $time);
            error();
        end
        @(posedge clk);
        #1step;
        if (RegWrite)
            regfile.write_reg_i(instruction, tb_writeData);
        if (PCSrc) tb_PC = tb_PC + cur_inst.imm_b();
        else tb_PC = tb_PC + 4;
        RegWrite = 0;
        loadPC = 0;
    endtask

    // Data path
    // assign PCSrc = tb_alu_Zero & riscv_ctrl.branch;
    // assign writeData = MemtoReg ? dReadData : tb_alu;

    initial begin
        regfile = new();
        inst_mem = new(MAX_TEXT_SIZE, instruction_memory_filename);
        data_mem = new(MAX_DATA_SIZE, data_memory_filename);

        //shall print %t with scaled in ns (-9), with 2 precision digits, and would print the " ns" string
        $timeformat(-9, 0, " ns", 20);
        $display("*** Start of Simulation ***");
        
        // Initialize the inputs
        repeat(3) @(negedge clk);
        rst = 0;
        repeat(3) @(negedge clk);
        // Default control signals
        init_control();

        // Issue a global reset
        rst = 1;
        tb_PC = TB_INITIAL_PC;
        repeat(3) @(negedge clk);
        rst = 0;
        repeat(3) @(negedge clk);

        init_control();
        
        repeat(3) @(negedge clk);

        @(posedge clk);
        while(instruction != riscv_instr::EBREAK_INSTRUCTION)
            execute_instruction();
        init_control();

        repeat(20) @(negedge clk);

        $display("*** Simulation done *** %0t", $time);
        $display("===== TEST PASSED =====");

        $finish;

    end  // end initial
    
endmodule